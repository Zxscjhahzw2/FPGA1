library verilog;
use verilog.vl_types.all;
entity rgy_vlg_vec_tst is
end rgy_vlg_vec_tst;
